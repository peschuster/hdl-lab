library verilog;
use verilog.vl_types.all;
entity decode_tb is
end decode_tb;
