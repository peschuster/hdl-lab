// Integrated Electronic Systems Lab
// TU Darmstadt
// Author:	Group 6
// Email:
//
// ALU Module.
// Computes add, sub, mv and cmp command
 // For cmp using the sub command code

// sel_in mapping
// using bit 1 to 3 of first byte 
// 000 - add
// 101 - sub
// 001 - mv (imm)
// 010 - mv (reg)

// apsr
// 31 30 29 28
// N  Z  C  V
// mapped to
// 3 2 1 0
// N Z C V
//
//N - 1 if result of rn - imm < 0; 0 else
//Z - 1 if result of rn - imm = 0; 0 else
// not implemented yet:
//C - 1 if results in a carry condition (unsigned overflow); 0 else
//V - 1 if results in a overflow condition (signed overflow); 0 else

module alu(
	i_imm,
	i_rn,
	i_sel,
	o_result,
	o_apsr
);

input logic [31:0] 	i_imm;
input logic [31:0] 	i_rn;
input logic [2:0]   i_sel;

output logic [31:0] 	o_result;
output logic [3:0]    o_apsr;

logic [32:0]  iresult_r; 


always@ (*) begin
  //reset APSR
  o_apsr = 0;

  //calculate
  case (i_sel)
    3'b000:
      //add
		  iresult_r = i_imm + i_rn;
    3'b101: begin
      //sub
		  iresult_r = i_rn - i_imm;
      if (iresult_r[32] == 1'b1) begin
        o_apsr[3] = 1;
      end
    end
    3'b001:
      //mv (imm)
      iresult_r = i_imm;
    3'b010:
      //mv (reg)
      iresult_r = i_rn;
    default:
      // error
      iresult_r = 0;
  endcase

  // set intermal result to output result
  o_result = iresult_r[31:0];

  if (o_result == 0) begin
    //set Z flag
    o_apsr[2] = 1;
  end
 
end

endmodule
