library verilog;
use verilog.vl_types.all;
entity ir_cache_ctrl_tb is
end ir_cache_ctrl_tb;
